`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   08:28:48 12/13/2019
// Design Name:   booth
// Module Name:   D:/Aanshi/AANSHI PATWARI-2019/Semester 3/booth_algorithm/booth_tb.v
// Project Name:  booth_algorithm
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: booth
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module booth_tb;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	booth uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

